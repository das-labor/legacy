-- DDR controller
  constant CFG_DDRSP  		: integer := CONFIG_DDRSP;
  constant CFG_DDRSP_INIT  	: integer := CONFIG_DDRSP_INIT;
  constant CFG_DDRSP_FREQ   	: integer := CONFIG_DDRSP_FREQ;
  constant CFG_DDRSP_COL    	: integer := CONFIG_DDRSP_COL;
  constant CFG_DDRSP_SIZE  	: integer := CONFIG_DDRSP_SIZE;

