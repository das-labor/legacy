library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;



entity f_eins is
    Port ( f1 : out  STD_LOGIC);
end f_eins;

architecture Behavioral of f_eins is

begin

f1<='1';

end Behavioral;

