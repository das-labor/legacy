-----------------------------------------------------------------------------
-- Wishbone Block Ram -------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity wb_bram is
   port (
      clk      : in  std_logic;
      reset    : in  std_logic;
      -- Wishbone bus
      wb_adr_i : in  std_logic_vector(31 downto 0);
      wb_dat_i : in  std_logic_vector(31 downto 0);
      wb_dat_o : out std_logic_vector(31 downto 0);
      wb_sel_i : in  std_logic_vector( 3 downto 0);
      wb_cyc_i : in  std_logic;
      wb_stb_i : in  std_logic;
      wb_ack_o : out std_logic;
      wb_we_i  : in  std_logic );
end wb_bram;

-----------------------------------------------------------------------------
-- Implementation -----------------------------------------------------------
architecture rtl of wb_bram is

constant mem_size : natural := (1*512) - 1;
type mem_type is array(0 to mem_size) of std_logic_vector(31 downto 0);

-----------------------------------------------------------------------------
-- Pre-Initialized-Data -----------------------------------------------------
signal mem : mem_type := (

     x"88100000", x"09000000", x"81c12200", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"91d02000", x"01000000", x"01000000", x"01000000", 
     x"ae102001", x"a1480000", x"1080004e", x"a7500000", 
     x"ae102002", x"a1480000", x"1080004a", x"a7500000", 
     x"ae102003", x"a1480000", x"10800046", x"a7500000", 
     x"ae102004", x"a1480000", x"10800042", x"a7500000", 
     x"ae102005", x"a1480000", x"1080003e", x"a7500000", 
     x"ae102006", x"a1480000", x"1080003a", x"a7500000", 
     x"ae102007", x"a1480000", x"10800036", x"a7500000", 
     x"ae102008", x"a1480000", x"10800032", x"a7500000", 
     x"ae102009", x"a1480000", x"1080002e", x"a7500000", 
     x"ae10200a", x"a1480000", x"1080002a", x"a7500000", 
     x"ae10200b", x"a1480000", x"10800026", x"a7500000", 
     x"ae10200c", x"a1480000", x"10800022", x"a7500000", 
     x"ae10200d", x"a1480000", x"1080001e", x"a7500000", 
     x"ae10200e", x"a1480000", x"1080001a", x"a7500000", 
     x"ae10200f", x"a1480000", x"10800016", x"a7500000", 
     x"821020c0", x"81884000", x"05000000", x"8410a000", 
     x"81988000", x"84006001", x"8408a007", x"86102001", 
     x"8728c002", x"8190c000", x"3d20ffff", x"bc17a3fc", 
     x"bc2fa00f", x"9c27a040", x"82106020", x"81884000", 
     x"92100000", x"90100000", x"40000050", x"01000000", 
     x"4000009d", x"90100017", x"81c44000", x"81cc8000", 
     x"a7800000", x"81c3e008", x"01000000", x"91480000", 
     x"902a2f00", x"81c3e008", x"818a0000", x"91480000", 
     x"90122f20", x"81c3e008", x"818a0000", x"81c20000", 
     x"01000000", x"9de3bf98", x"400000ef", x"01000000", 
     x"400000ed", x"b00a20ff", x"900a20ff", x"b12e2008", 
     x"400000e9", x"b0060008", x"900a20ff", x"b12e2008", 
     x"400000e5", x"b0060008", x"900a20ff", x"b12e2008", 
     x"81c7e008", x"91ee0008", x"9de3bf98", x"233c0000", 
     x"a0102007", x"920e0011", x"9332601c", x"90026030", 
     x"80a26009", x"04800003", x"94026037", x"9010000a", 
     x"400000f9", x"b12e2004", x"a0843fff", x"1cbffff7", 
     x"920e0011", x"01000000", x"81c7e008", x"81e80000", 
     x"9de3bf98", x"1120003f", x"901223fe", x"21200000", 
     x"e0240000", x"a0042004", x"80a40008", x"28bffffe", 
     x"e0240000", x"1120003f", x"a41223fe", x"21200000", 
     x"23000001", x"d2040000", x"901463a0", x"80a24010", 
     x"02800004", x"a0042004", x"400000f9", x"01000000", 
     x"80a40012", x"28bffff9", x"d2040000", x"01000000", 
     x"81c7e008", x"81e80000", x"9de3bf98", x"133c0400", 
     x"90102023", x"92126010", x"4000009f", x"d02a4000", 
     x"7fffffb3", x"01000000", x"11000001", x"400000e8", 
     x"901223b8", x"7fffffdb", x"01000000", x"400000a6", 
     x"01000000", x"912a2018", x"913a2018", x"80a22072", 
     x"02800038", x"01000000", x"04800024", x"80a22075", 
     x"12bffff7", x"11000001", x"400000d9", x"901223d8", 
     x"7fffffa9", x"01000000", x"7fffffb8", x"a2100008", 
     x"400000b9", x"9010203a", x"7fffffa3", x"01000000", 
     x"7fffffb2", x"a0100008", x"9010203a", x"400000b2", 
     x"a4044010", x"80a44012", x"1a80000a", x"a0102000", 
     x"40000089", x"01000000", x"d02c4000", x"900a20ff", 
     x"a2046001", x"80a44012", x"0abffffa", x"a0040008", 
     x"7fffffa2", x"90100010", x"11000001", x"901223e0", 
     x"400000bb", x"9e03ff54", x"80a22067", x"12bfffd4", 
     x"11000001", x"400000b6", x"901223e8", x"7fffff86", 
     x"01000000", x"7fffff95", x"a2100008", x"40000096", 
     x"9010202e", x"7fffff7a", x"01000000", x"7fffff7c", 
     x"90100011", x"11000001", x"10bfffee", x"901223f0", 
     x"7fffff77", x"90102000", x"10bfffcc", x"11000001", 
     x"01000000", x"80a22006", x"0280002a", x"01000000", 
     x"08800028", x"80a2200a", x"0280000b", x"80a2200c", 
     x"12800024", x"11000001", x"d4022398", x"13000001", 
     x"d002639c", x"d6028000", x"90022001", x"1080001d", 
     x"d022639c", x"1920c000", x"d4032020", x"1320c000", 
     x"d0026024", x"94a28008", x"2c800002", x"9402a020", 
     x"80a2a01e", x"14800011", x"11000001", x"d6032020", 
     x"d4022394", x"d202a008", x"d22ac000", x"d0032020", 
     x"90022001", x"d0232020", x"d2032020", x"1120c000", 
     x"90122020", x"80a24008", x"12800006", x"90027fe0", 
     x"d0232020", x"30800003", x"d2022394", x"d4026008", 
     x"01000000", x"81c3e008", x"01000000", x"9de3bf98", 
     x"912e2001", x"90020018", x"932a2006", x"90020009", 
     x"912a2002", x"90020018", x"15000001", x"912a2002", 
     x"d202a398", x"90020018", x"912a2004", x"d0226010", 
     x"c0226014", x"9010200a", x"d022600c", x"b010000a", 
     x"7fffff28", x"01000000", x"d0062398", x"d202200c", 
     x"808a6001", x"02bffffb", x"01000000", x"01000000", 
     x"81c7e008", x"81e80000", x"13000001", x"d4026398", 
     x"11000030", x"90122350", x"d022a004", x"c022a008", 
     x"9010200e", x"d0228000", x"01000000", x"81c3e008", 
     x"01000000", x"11000001", x"d8022394", x"921021b2", 
     x"1120c000", x"d2232004", x"1720c000", x"90122000", 
     x"d022e024", x"d402e024", x"1120c000", x"d4222020", 
     x"92102004", x"d2230000", x"01000000", x"81c3e008", 
     x"01000000", x"9de3bf98", x"1720c000", x"d202e020", 
     x"1520c000", x"d002a024", x"80a24008", x"02800011", 
     x"a010000b", x"d002a024", x"f00a0000", x"d202a024", 
     x"1120c000", x"92026001", x"d222a024", x"d202a024", 
     x"90122020", x"80a24008", x"3280000f", x"b12e2018", 
     x"90027fe0", x"d022a024", x"1080000b", x"b12e2018", 
     x"b010000a", x"7ffffeeb", x"01000000", x"d2042020", 
     x"d0062024", x"80a24008", x"02bffffb", x"1520c000", 
     x"30bfffe9", x"b13e2018", x"01000000", x"81c7e008", 
     x"81e80000", x"9de3bf98", x"23000001", x"d2046394", 
     x"d0024000", x"808a2002", x"2280000c", x"13000001", 
     x"a010200c", x"e0224000", x"7ffffed6", x"01000000", 
     x"d2046394", x"d0024000", x"808a2002", x"12bffffa", 
     x"01000000", x"13000001", x"d4026394", x"912e2018", 
     x"913a2018", x"d022a008", x"92102004", x"d2228000", 
     x"01000000", x"81c7e008", x"81e80000", x"9de3bf98", 
     x"d00e0000", x"912a2018", x"80a22000", x"0280000a", 
     x"01000000", x"7fffffe0", x"913a2018", x"b0062001", 
     x"d00e0000", x"912a2018", x"80a22000", x"12bffffa", 
     x"01000000", x"01000000", x"81c7e008", x"81e80000", 
     x"f0000000", x"f0010000", x"f0020000", x"00000000", 
     x"44445220", x"54455354", x"20464149", x"4c45440a", 
     x"00000000", x"00000000", x"0d0a2a2a", x"20535049", 
     x"4b452042", x"4f4f544c", x"4f414445", x"52202a2a", 
     x"0a0d0000", x"00000000", x"753a0000", x"00000000", 
     x"2e0d0a00", x"00000000", x"673a0000", x"00000000", 
     x"58585858", x"00000000", 


    others => x"00000000" 
);
	
signal ack : std_logic;

begin

wb_ack_o <= wb_stb_i and ack;

memproc: process (clk) is
variable a : integer;
begin
	if clk'event and clk='1' then
	if wb_stb_i='1' then
		a := to_integer(unsigned(wb_adr_i(15 downto 2)));
	
		if wb_we_i='1' then 
			mem(a) <= wb_dat_i;
		end if;
		
--			if wb_sel_i(3)='1' then
--				mem(a)(31 downto 24) <= wb_dat_i(31 downto 24);
--			end if;
--			if wb_sel_i(2)='1' then
--				mem(a)(23 downto 16) <= wb_dat_i(23 downto 16);
--			end if;
--			if wb_sel_i(1)='1' then
--				mem(a)(15 downto  8) <= wb_dat_i(15 downto  8);
--			end if;
--			if wb_sel_i(0)='1' then
--				mem(a)( 7 downto  0) <= wb_dat_i( 7 downto  0);
--			end if;
--		end if;


		wb_dat_o <= mem(a);
		ack <= '1' and not ack;
	else
		ack <= '0';
	end if;
	end if;
end process;

end rtl;

