-- USB target controller
  constant CFG_USBDCL     	: integer := CONFIG_USBDCL;

