-- ATA interface
  constant CFG_ATA      : integer := CONFIG_ATA_ENABLE;
  constant CFG_ATAIO    : integer := 16#CONFIG_ATAIO#;
  constant CFG_ATAIRQ   : integer := CONFIG_ATAIRQ;

