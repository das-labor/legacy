-- pragma translate_off
use std.textio.all;
-- pragma translate_on
package version is
  constant grlib_version : integer := 1010;
-- pragma translate_off
  constant grlib_date : string := "20060909";
-- pragma translate_on
  constant grlib_build : integer := 1640;
end;
