
library ieee;
use ieee.std_logic_1164.all;

use ieee.numeric_std.all;

entity rom is
port (addr	:in std_logic_vector (10 downto 0);
        data  :out std_logic_vector (15 downto 0); 
		clk  : in std_logic		);
end rom;


architecture rtl of rom is
	type rom_array is array (0 to 2047) of std_logic_vector(15 downto 0);
constant ROM : ROM_ARRAY := (
		x"94F8",x"EF8F",x"E09F",x"BF8D",x"BF9E",x"940E",x"F8B5",x"940E"
		,x"F8E4",x"2799",x"368D",x"0591",x"F409",x"C077",x"368E",x"0591"
		,x"F484",x"3684",x"0591",x"F409",x"C055",x"3685",x"0591",x"F424"
		,x"3682",x"0591",x"F1C1",x"CFEB",x"368A",x"0591",x"F409",x"C08C"
		,x"CFE6",x"3784",x"0591",x"F409",x"C07D",x"3785",x"0591",x"F42C"
		,x"3782",x"0591",x"F409",x"C085",x"CFDA",x"3785",x"0591",x"F6B9"
		,x"940E",x"F8F8",x"2F08",x"2F19",x"940E",x"F8F8",x"2FD9",x"2FC8"
		,x"9721",x"EF8F",x"3FCF",x"07D8",x"F251",x"2F81",x"2799",x"5080"
		,x"4F9E",x"9390",x"FE01",x"9380",x"FE00",x"940E",x"F8E4",x"2FF1"
		,x"2FE0",x"6FFF",x"8380",x"5F0F",x"4F1F",x"9721",x"EFEF",x"3FCF"
		,x"07DE",x"F759",x"CFB4",x"940E",x"F8F8",x"2F08",x"2F19",x"940E"
		,x"F8F8",x"2FD9",x"2FC8",x"9721",x"EFFF",x"3FCF",x"07DF",x"F409"
		,x"CFA6",x"2FF1",x"2FE0",x"95C8",x"2D80",x"940E",x"F8BA",x"5F0F"
		,x"4F1F",x"CFF1",x"940E",x"F8F8",x"2F08",x"2F19",x"940E",x"F8F8"
		,x"2FD9",x"2FC8",x"9721",x"EF8F",x"3FCF",x"07D8",x"F409",x"CF8F"
		,x"2FF1",x"2FE0",x"9181",x"2F0E",x"2F1F",x"940E",x"F8BA",x"9721"
		,x"EFFF",x"3FCF",x"07DF",x"F7A1",x"CF82",x"E0C0",x"EF8F",x"2FEC"
		,x"27FF",x"50E0",x"47F0",x"93C1",x"8380",x"5FCE",x"3FCE",x"F7B9"
		,x"E0C0",x"2FEC",x"27FF",x"50E0",x"47F0",x"8180",x"178C",x"F031"
		,x"E686",x"940E",x"F8BA",x"2F8C",x"940E",x"F8BA",x"5FCE",x"3FCE"
		,x"F781",x"CF65",x"E0C0",x"E0D0",x"2F8C",x"940E",x"F8BA",x"9621"
		,x"3FCF",x"05D1",x"F3C9",x"F3C0",x"940E",x"F8F8",x"2FE8",x"2FF9"
		,x"9509",x"E782",x"940E",x"F8BA",x"CF52",x"9A53",x"9A54",x"E188"
		,x"B989",x"9508",x"9B5D",x"CFFE",x"B98C",x"9508",x"93CF",x"93DF"
		,x"2FD9",x"2FC8",x"8188",x"2388",x"F031",x"9189",x"940E",x"F8BA"
		,x"8188",x"2388",x"F7D1",x"91DF",x"91CF",x"9508",x"93CF",x"93DF"
		,x"2FD9",x"2FC8",x"2FF9",x"2FE8",x"95C8",x"2D80",x"2388",x"F049"
		,x"940E",x"F8BA",x"9621",x"2FFD",x"2FEC",x"95C8",x"2D80",x"2388"
		,x"F7B9",x"91DF",x"91CF",x"9508",x"9B5F",x"CFFE",x"B18C",x"2799"
		,x"FD87",x"9590",x"9508",x"2FF9",x"2FE8",x"9B5F",x"C005",x"B18C"
		,x"8380",x"E081",x"E090",x"9508",x"E080",x"E090",x"9508",x"9508"
		,x"930F",x"931F",x"940E",x"F8E4",x"2F08",x"940E",x"F8E4",x"2F18"
		,x"2F91",x"2F80",x"911F",x"910F",x"9508",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
		,x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000"
			);
begin
	p_rom : process(clk, addr)
	begin
	if clk'event and clk = '0' then
		data <= ROM(to_integer(unsigned(addr)));
	end if;
	end process;
end rtl;
