-- MIL-STD-1553 controllers

  constant CFG_1553_RT_EN         : integer := CONFIG_1553_RT_EN;
  constant CFG_1553_RTADDR        : integer := CONFIG_1553_RTADDR;
  constant CFG_1553_RTADDRP    	  : integer := CONFIG_1553_RTADDRP;
  constant CFG_1553_WRTCMD    	  : integer := CONFIG_1553_WRTCMD;
  constant CFG_1553_WRTTSW        : integer := CONFIG_1553_WRTTSW;
  constant CFG_1553_INTENBBR      : integer := CONFIG_1553_INTENBBR;
  constant CFG_1553_BCASTEN    	  : integer := CONFIG_1553_BCASTEN;
  constant CFG_1553_SA30LOOP      : integer := CONFIG_1553_SA30LOOP;
  constant CFG_1553_RTCLKSPD      : integer :=CONFIG_1553_RTCLKSPD;
  constant CFG_1553_BC_EN         : integer := CONFIG_1553_BC_EN;
  constant CFG_1553_BRM_EN        : integer := CONFIG_1553_BRM_EN;
  constant CFG_1553_NUM           : integer := CONFIG_1553_NUM;
  constant CFG_1553_BRM_ABSTD     : integer := CONFIG_1553_BRM_ABSTD;
  constant CFG_1553_BRM_MS    	  : integer := CONFIG_1553_BRM_MS;

  
