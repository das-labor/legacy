-- Gaisler Ethernet core
  constant CFG_GRETH   	: integer := CONFIG_GRETH_ENABLE;
  constant CFG_ETH_FIFO : integer := CFG_GRETH_FIFO;

