-----------------------------------------------------------------------------
-- Wishbone Block Ram -------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity wb_bram is
   port (
      clk      : in  std_logic;
      reset    : in  std_logic;
      -- Wishbone bus
      wb_adr_i : in  std_logic_vector(31 downto 0);
      wb_dat_i : in  std_logic_vector(31 downto 0);
      wb_dat_o : out std_logic_vector(31 downto 0);
      wb_sel_i : in  std_logic_vector( 3 downto 0);
      wb_cyc_i : in  std_logic;
      wb_stb_i : in  std_logic;
      wb_ack_o : out std_logic;
      wb_we_i  : in  std_logic );
end wb_bram;

-----------------------------------------------------------------------------
-- Implementation -----------------------------------------------------------
architecture rtl of wb_bram is

constant mem_size : natural := (8*512) - 1;
type mem_type is array(0 to mem_size) of std_logic_vector(31 downto 0);

-----------------------------------------------------------------------------
-- Pre-Initialized-Data -----------------------------------------------------
signal mem : mem_type := (
     x"98000000", x"d0000000", x"78010000", x"38210000", 
     x"d0e10000", x"f8000003", x"34000000", x"34000000", 
     x"98000000", x"781c0000", x"3b9c1000", x"379cfffc", 
     x"781a0000", x"3b5a0800", x"34010000", x"34020000", 
     x"34030000", x"f800006f", x"c3a00000", x"c3a00000", 
     x"e0000000", x"e0000000", x"379cff80", x"5b810004", 
     x"5b820008", x"5b83000c", x"5b840010", x"5b850014", 
     x"5b860018", x"5b87001c", x"5b880020", x"5b890024", 
     x"5b8a0028", x"5b9e0078", x"5b9f007c", x"2b810080", 
     x"5b810074", x"bb800800", x"34210080", x"5b810070", 
     x"c3a00000", x"2b810004", x"2b820008", x"2b83000c", 
     x"2b840010", x"2b850014", x"2b860018", x"2b87001c", 
     x"2b880020", x"2b890024", x"2b8a0028", x"2b9d0074", 
     x"2b9e0078", x"2b9f007c", x"2b9c0070", x"c3c00000", 
     x"379cfff8", x"5b8b0008", x"5b9d0004", x"f80000ee", 
     x"3c2b0008", x"f80000ec", x"b5615800", x"3d6b0008", 
     x"f80000e9", x"b5615800", x"3d6b0008", x"f80000e6", 
     x"b5610800", x"2b8b0008", x"2b9d0004", x"379c0008", 
     x"c3a00000", x"379cfff0", x"5b8b0010", x"5b8c000c", 
     x"5b8d0008", x"5b9d0004", x"780df000", x"b8205800", 
     x"39ad0000", x"340c0007", x"a16d0800", x"0023001c", 
     x"68620009", x"34610030", x"44400002", x"34610037", 
     x"3d6b0004", x"f8000101", x"358cffff", x"4d80fff7", 
     x"2b8b0010", x"2b8c000c", x"2b8d0008", x"2b9d0004", 
     x"379c0010", x"c3a00000", x"379cfff4", x"5b8b000c", 
     x"5b8c0008", x"5b9d0004", x"780b8000", x"b9601000", 
     x"78018000", x"396b0000", x"3821fffe", x"596b0000", 
     x"356b0004", x"55610002", x"e3fffffd", x"b8405800", 
     x"780c8000", x"396b0000", x"398cfffe", x"29620000", 
     x"78010000", x"38210638", x"444b0002", x"f8000106", 
     x"356b0004", x"556c0002", x"e3fffff9", x"2b8b000c", 
     x"2b8c0008", x"2b9d0004", x"379c000c", x"c3a00000", 
     x"379cffec", x"5b8b0014", x"5b8c0010", x"5b8d000c", 
     x"5b8e0008", x"5b9d0004", x"f8000092", x"fbffff8b", 
     x"78010000", x"3821064c", x"f80000f3", x"fbffffd7", 
     x"f800009d", x"b8201000", x"64210072", x"5c200017", 
     x"68410072", x"5c20002e", x"64410067", x"4420fff9", 
     x"78010000", x"38210668", x"f80000e7", x"fbffffa1", 
     x"b8207000", x"fbffffb0", x"3401002e", x"f80000bf", 
     x"fbffff77", x"b9c00800", x"fbffff76", x"78010000", 
     x"3821066c", x"f80000dc", x"f8000087", x"b8201000", 
     x"64210072", x"4420ffeb", x"34010000", x"fbffff6d", 
     x"78010000", x"38210674", x"f80000d3", x"fbffff8d", 
     x"b8207000", x"fbffff9c", x"3401003a", x"f80000ab", 
     x"fbffff88", x"b8205800", x"fbffff97", x"3401003a", 
     x"b5cb6800", x"f80000a5", x"340c0000", x"b9c05800", 
     x"51cd000a", x"f8000070", x"31610000", x"b5816000", 
     x"356b0001", x"516d0005", x"e3fffffb", x"64410075", 
     x"4420ffcc", x"e3ffffe7", x"b9800800", x"fbffff86", 
     x"78010000", x"38210678", x"f80000b7", x"e3ffffdb", 
     x"6422000c", x"78040000", x"78030000", x"6421000a", 
     x"38840820", x"38630824", x"5c20000d", x"78010000", 
     x"78040000", x"38210634", x"38840628", x"5c400002", 
     x"c3a00000", x"28210000", x"28820000", x"28230000", 
     x"34420001", x"58820000", x"c3a00000", x"28820000", 
     x"78060000", x"38c60630", x"28610000", x"78070000", 
     x"b8c02800", x"38e70820", x"c8410800", x"4c200002", 
     x"34210020", x"6821001e", x"5c20000e", x"28830000", 
     x"28c10000", x"78050000", x"38a50800", x"28220008", 
     x"30620000", x"28810000", x"34210001", x"58810000", 
     x"28820000", x"5c47ffe3", x"58850000", x"c3a00000", 
     x"28a10000", x"28220008", x"c3a00000", x"379cfff8", 
     x"5b8b0008", x"5b9d0004", x"78040000", x"38840634", 
     x"3802c350", x"88220800", x"28830000", x"b8805800", 
     x"3402000a", x"58610010", x"34010000", x"58610014", 
     x"5862000c", x"fbffff10", x"29620000", x"2841000c", 
     x"20210001", x"4420fffc", x"2b8b0008", x"2b9d0004", 
     x"379c0008", x"c3a00000", x"78010000", x"38210634", 
     x"28230000", x"3802c350", x"58620004", x"34010000", 
     x"58610008", x"3402000e", x"58620000", x"c3a00000", 
     x"78010000", x"38210630", x"28250000", x"78030000", 
     x"78020000", x"340101b2", x"58a10004", x"38630824", 
     x"38420800", x"58620000", x"28640000", x"78010000", 
     x"38210820", x"58240000", x"34020004", x"58a20000", 
     x"c3a00000", x"379cfff0", x"5b8b0010", x"5b8c000c", 
     x"5b8d0008", x"5b9d0004", x"78030000", x"38630820", 
     x"28620000", x"780d0000", x"b9a02000", x"38840824", 
     x"28810000", x"44410014", x"b9a02800", x"38a50824", 
     x"28a40000", x"78030000", x"38630820", x"40820000", 
     x"28a10000", x"204400ff", x"34210001", x"58a10000", 
     x"28a20000", x"4443000f", x"b8800800", x"2b8b0010", 
     x"2b8c000c", x"2b8d0008", x"2b9d0004", x"379c0010", 
     x"c3a00000", x"b8606000", x"b8805800", x"fbfffeca", 
     x"29820000", x"29610000", x"4441fffd", x"e3ffffe7", 
     x"78010000", x"38210800", x"58a10000", x"b8800800", 
     x"2b8b0010", x"2b8c000c", x"2b8d0008", x"2b9d0004", 
     x"379c0010", x"c3a00000", x"379cffec", x"5b8b0014", 
     x"5b8c0010", x"5b8d000c", x"5b8e0008", x"5b9d0004", 
     x"780d0000", x"b9a01800", x"38630630", x"28620000", 
     x"202e00ff", x"28410000", x"20210002", x"4420000a", 
     x"b8605800", x"340c000c", x"29610000", x"582c0000", 
     x"fbfffea9", x"29620000", x"28410000", x"20210002", 
     x"5c20fffa", x"39ad0630", x"29a20000", x"34010004", 
     x"584e0008", x"58410000", x"2b8b0014", x"2b8c0010", 
     x"2b8d000c", x"2b8e0008", x"2b9d0004", x"379c0014", 
     x"c3a00000", x"379cfff8", x"5b8b0008", x"5b9d0004", 
     x"b8205800", x"e0000003", x"fbffffd8", x"356b0001", 
     x"41610000", x"5c20fffd", x"2b8b0008", x"2b9d0004", 
     x"379c0008", x"c3a00000", x"00000000", x"80002000", 
     x"80001000", x"80000000", x"44445220", x"54455354", 
     x"20464149", x"4c45440a", x"00000000", x"0d0a2a2a", 
     x"20535049", x"4b452042", x"4f4f544c", x"4f414445", 
     x"52202a2a", x"0a0d0000", x"673a0000", x"58585858", 
     x"00000000", x"753a0000", x"2e0d0a00", 


   others => x"00000000" 
);
	
signal ack : std_logic;

begin

wb_ack_o <= wb_stb_i and ack;

memproc: process (clk) is
variable a : integer;
begin
	if clk'event and clk='1' then
	if wb_stb_i='1' and wb_cyc_i='1' then
		a := to_integer(unsigned(wb_adr_i(12 downto 2)));
	
		if wb_we_i='1' then 
			mem(a) <= wb_dat_i;
		end if;
		
--			if wb_sel_i(3)='1' then
--				mem(a)(31 downto 24) <= wb_dat_i(31 downto 24);
--			end if;
--			if wb_sel_i(2)='1' then
--				mem(a)(23 downto 16) <= wb_dat_i(23 downto 16);
--			end if;
--			if wb_sel_i(1)='1' then
--				mem(a)(15 downto  8) <= wb_dat_i(15 downto  8);
--			end if;
--			if wb_sel_i(0)='1' then
--				mem(a)( 7 downto  0) <= wb_dat_i( 7 downto  0);
--			end if;
--		end if;


		wb_dat_o <= mem(a);
		ack <= '1' and not ack after 2 ns;
	else
		ack <= '0';
	end if;
	end if;
end process;

end rtl;

