-- LEON2 memory controller
  constant CFG_MCTRL_LEON2    : integer := CONFIG_MCTRL_LEON2;
  constant CFG_MCTRL_RAM8BIT  : integer := CONFIG_MCTRL_8BIT;
  constant CFG_MCTRL_RAM16BIT : integer := CONFIG_MCTRL_16BIT;
  constant CFG_MCTRL_5CS      : integer := CONFIG_MCTRL_5CS;
  constant CFG_MCTRL_SDEN    	: integer := CONFIG_MCTRL_SDRAM;
  constant CFG_MCTRL_SEPBUS  	: integer := CONFIG_MCTRL_SDRAM_SEPBUS;
  constant CFG_MCTRL_INVCLK  	: integer := CONFIG_MCTRL_SDRAM_INVCLK;
  constant CFG_MCTRL_SD64    	: integer := CONFIG_MCTRL_SDRAM_BUS64;

