-- SSRAM controller
  constant CFG_SSCTRL  	: integer := CONFIG_SSCTRL;

