-- VGA and PS2/ interface
  constant CFG_KBD_ENABLE : integer := CONFIG_KBD_ENABLE;
  constant CFG_VGA_ENABLE : integer := CONFIG_VGA_ENABLE;

