-- PROM/SRAM controller
  constant CFG_SRCTRL         	: integer := CONFIG_SRCTRL;
  constant CFG_SRCTRL_PROMWS  	: integer := CONFIG_SRCTRL_PROMWS;
  constant CFG_SRCTRL_RAMWS   	: integer := CONFIG_SRCTRL_RAMWS;
  constant CFG_SRCTRL_RMW  	: integer := CONFIG_SRCTRL_RMW;
  constant CFG_SRCTRL_8BIT    	: integer := CONFIG_SRCTRL_8BIT;

