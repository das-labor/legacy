-- USB target controller
  constant CFG_USBTGT     	: integer := CONFIG_USBTGT;

