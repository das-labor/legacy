-- AMBA settings
  constant CFG_DEFMST  	: integer := CONFIG_AHB_DEFMST;
  constant CFG_RROBIN  	: integer := CONFIG_AHB_RROBIN;
  constant CFG_SPLIT   	: integer := CONFIG_AHB_SPLIT;
  constant CFG_AHBIO   	: integer := 16#CONFIG_AHB_IOADDR#;
  constant CFG_APBADDR 	: integer := 16#CONFIG_APB_HADDR#;

